`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:28:03 10/09/2017 
// Design Name: 
// Module Name:    DEMUX1_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DEMUX1_2(
    input [7:0] Data_in,
    input Select_line,
    input CLK,
    input RESET,
    output [7:0] OUT_A,
    output [7:0] OUT_B
    );


endmodule
